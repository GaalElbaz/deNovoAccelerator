module topDesgin_tbFive();

	logic clk, rstN;
	logic [31:0] randA;
	logic [31:0] randB;
	logic unsigned [48:0][31:0] kmersSeqOne;
	logic unsigned [48:0][31:0] kmersSeqTwo;
	logic unsigned [4:0] jaccardSimilarity;
	
	topDesginModule myTopDesginTB(.clk(clk), .rstN(rstN), .randA(randA), .randB(randB), .kmersSeqOne(kmersSeqOne), .kmersSeqTwo(kmersSeqTwo), .jaccardSimilarity(jaccardSimilarity));
	
	always begin
		#40 clk = ~clk;
	end
	
	initial begin
		clk = 0;
		rstN = 1;
		kmersSeqOne[0]= 32'b11000110100011111000111100100001;
		kmersSeqOne[1]= 32'b00011010001111100011110010000111;
		kmersSeqOne[2]= 32'b01101000111110001111001000011100;
		kmersSeqOne[3]= 32'b10100011111000111100100001110001;
		kmersSeqOne[4]= 32'b10001111100011110010000111000110;
		kmersSeqOne[5]= 32'b00111110001111001000011100011010;
		kmersSeqOne[6]= 32'b11111000111100100001110001101000;
		kmersSeqOne[7]= 32'b11100011110010000111000110100011;
		kmersSeqOne[8]= 32'b10001111001000011100011010001111;
		kmersSeqOne[9]= 32'b00111100100001110001101000111110;
		kmersSeqOne[10]= 32'b11110010000111000110100011111000;
		kmersSeqOne[11]= 32'b11001000011100011010001111100011;
		kmersSeqOne[12]= 32'b00100001110001101000111110001111;
		kmersSeqOne[13]= 32'b10000111000110100011111000111100;
		kmersSeqOne[14]= 32'b00011100011010001111100011110010;
		kmersSeqOne[15]= 32'b01110001101000111110001111001000;
		kmersSeqOne[16]= 32'b11000110100011111000111100100001;
		kmersSeqOne[17]= 32'b00011010001111100011110010000110;
		kmersSeqOne[18]= 32'b01101000111110001111001000011011;
		kmersSeqOne[19]= 32'b10100011111000111100100001101100;
		kmersSeqOne[20]= 32'b10001111100011110010000110110010;
		kmersSeqOne[21]= 32'b00111110001111001000011011001001;
		kmersSeqOne[22]= 32'b11111000111100100001101100100100;
		kmersSeqOne[23]= 32'b11100011110010000110110010010011;
		kmersSeqOne[24]= 32'b10001111001000011011001001001111;
		kmersSeqOne[25]= 32'b00111100100001101100100100111110;
		kmersSeqOne[26]= 32'b11110010000110110010010011111000;
		kmersSeqOne[27]= 32'b11001000011011001001001111100011;
		kmersSeqOne[28]= 32'b00100001101100100100111110001111;
		kmersSeqOne[29]= 32'b10000110110010010011111000111100;
		kmersSeqOne[30]= 32'b00011011001001001111100011110010;
		kmersSeqOne[31]= 32'b01101100100100111110001111001000;
		kmersSeqOne[32]= 32'b10110010010011111000111100100001;
		kmersSeqOne[33]= 32'b11001001001111100011110010000101;
		kmersSeqOne[34]= 32'b00100100111110001111001000010110;
		kmersSeqOne[35]= 32'b10010011111000111100100001011001;
		kmersSeqOne[36]= 32'b01001111100011110010000101100110;
		kmersSeqOne[37]= 32'b00111110001111001000010110011001;
		kmersSeqOne[38]= 32'b11111000111100100001011001100110;
		kmersSeqOne[39]= 32'b11100011110010000101100110011001;
		kmersSeqOne[40]= 32'b10001111001000010110011001100110;
		kmersSeqOne[41]= 32'b00111100100001011001100110011001;
		kmersSeqOne[42]= 32'b11110010000101100110011001100110;
		kmersSeqOne[43]= 32'b11001000010110011001100110011001;
		kmersSeqOne[44]= 32'b00100001011001100110011001100110;
		kmersSeqOne[45]= 32'b10000101100110011001100110011001;
		kmersSeqOne[46]= 32'b00010110011001100110011001100110;
		kmersSeqOne[47]= 32'b01011001100110011001100110011001;
		kmersSeqOne[48]= 32'b01100110011001100110011001100110;
		kmersSeqTwo[0]= 32'b11000110100011111000011110010001;
		kmersSeqTwo[1]= 32'b00011010001111100001111001000110;
		kmersSeqTwo[2]= 32'b01101000111110000111100100011011;
		kmersSeqTwo[3]= 32'b10100011111000011110010001101100;
		kmersSeqTwo[4]= 32'b10001111100001111001000110110010;
		kmersSeqTwo[5]= 32'b00111110000111100100011011001010;
		kmersSeqTwo[6]= 32'b11111000011110010001101100101000;
		kmersSeqTwo[7]= 32'b11100001111001000110110010100011;
		kmersSeqTwo[8]= 32'b10000111100100011011001010001111;
		kmersSeqTwo[9]= 32'b00011110010001101100101000111110;
		kmersSeqTwo[10]= 32'b01111001000110110010100011111000;
		kmersSeqTwo[11]= 32'b11100100011011001010001111100001;
		kmersSeqTwo[12]= 32'b10010001101100101000111110000111;
		kmersSeqTwo[13]= 32'b01000110110010100011111000011110;
		kmersSeqTwo[14]= 32'b00011011001010001111100001111001;
		kmersSeqTwo[15]= 32'b01101100101000111110000111100100;
		kmersSeqTwo[16]= 32'b10110010100011111000011110010001;
		kmersSeqTwo[17]= 32'b11001010001111100001111001000110;
		kmersSeqTwo[18]= 32'b00101000111110000111100100011011;
		kmersSeqTwo[19]= 32'b10100011111000011110010001101100;
		kmersSeqTwo[20]= 32'b10001111100001111001000110110010;
		kmersSeqTwo[21]= 32'b00111110000111100100011011001001;
		kmersSeqTwo[22]= 32'b11111000011110010001101100100100;
		kmersSeqTwo[23]= 32'b11100001111001000110110010010011;
		kmersSeqTwo[24]= 32'b10000111100100011011001001001111;
		kmersSeqTwo[25]= 32'b00011110010001101100100100111110;
		kmersSeqTwo[26]= 32'b01111001000110110010010011111000;
		kmersSeqTwo[27]= 32'b11100100011011001001001111100001;
		kmersSeqTwo[28]= 32'b10010001101100100100111110000111;
		kmersSeqTwo[29]= 32'b01000110110010010011111000011110;
		kmersSeqTwo[30]= 32'b00011011001001001111100001111001;
		kmersSeqTwo[31]= 32'b01101100100100111110000111100100;
		kmersSeqTwo[32]= 32'b10110010010011111000011110010001;
		kmersSeqTwo[33]= 32'b11001001001111100001111001000101;
		kmersSeqTwo[34]= 32'b00100100111110000111100100010110;
		kmersSeqTwo[35]= 32'b10010011111000011110010001011001;
		kmersSeqTwo[36]= 32'b01001111100001111001000101100110;
		kmersSeqTwo[37]= 32'b00111110000111100100010110011001;
		kmersSeqTwo[38]= 32'b11111000011110010001011001100110;
		kmersSeqTwo[39]= 32'b11100001111001000101100110011001;
		kmersSeqTwo[40]= 32'b10000111100100010110011001100110;
		kmersSeqTwo[41]= 32'b00011110010001011001100110011001;
		kmersSeqTwo[42]= 32'b01111001000101100110011001100110;
		kmersSeqTwo[43]= 32'b11100100010110011001100110011001;
		kmersSeqTwo[44]= 32'b10010001011001100110011001100110;
		kmersSeqTwo[45]= 32'b01000101100110011001100110011001;
		kmersSeqTwo[46]= 32'b00010110011001100110011001100110;
		kmersSeqTwo[47]= 32'b01011001100110011001100110011001;
		kmersSeqTwo[48]= 32'b01100110011001100110011001100110;
		#20 rstN = 0;
		randA =  10323 ;
		randB =  10091 ;
		#80
		randA =  2324 ;
		randB =  1 ;
		#80
		randA =  358771 ;
		randB =  233 ;
		#80
		randA =  409712 ;
		randB =  76423 ;
		#80
		randA =  94390 ;
		randB =  4232409 ;
		#80
		randA =  2229481 ;
		randB =  57554 ;
		#80
		randA =  123 ;
		randB =  2231130 ;
		#80
		randA =  1441 ;
		randB =  1091 ;
		#260
		rstN = 1;
		$stop;
		$finish;
	end
	
	
	
	endmodule
	