module topDesgin_tbSix();

	logic clk, rstN;
	logic [31:0] randA;
	logic [31:0] randB;
	logic unsigned [48:0][31:0] kmersSeqOne;
	logic unsigned [48:0][31:0] kmersSeqTwo;
	logic unsigned [4:0] jaccardSimilarity;
	
	topDesginModule myTopDesginTB(.clk(clk), .rstN(rstN), .randA(randA), .randB(randB), .kmersSeqOne(kmersSeqOne), .kmersSeqTwo(kmersSeqTwo), .jaccardSimilarity(jaccardSimilarity));
	
	always begin
		#40 clk = ~clk;
	end
	
	initial begin
		clk = 0;
		rstN = 1;
		kmersSeqOne[0]= 32'b10000111101000010110111101001001;
		kmersSeqOne[1]= 32'b00011110100001011011110100100110;
		kmersSeqOne[2]= 32'b01111010000101101111010010011000;
		kmersSeqOne[3]= 32'b11101000010110111101001001100001;
		kmersSeqOne[4]= 32'b10100001011011110100100110000100;
		kmersSeqOne[5]= 32'b10000101101111010010011000010000;
		kmersSeqOne[6]= 32'b00010110111101001001100001000010;
		kmersSeqOne[7]= 32'b01011011110100100110000100001001;
		kmersSeqOne[8]= 32'b01101111010010011000010000100111;
		kmersSeqOne[9]= 32'b10111101001001100001000010011110;
		kmersSeqOne[10]= 32'b11110100100110000100001001111000;
		kmersSeqOne[11]= 32'b11010010011000010000100111100001;
		kmersSeqOne[12]= 32'b01001001100001000010011110000110;
		kmersSeqOne[13]= 32'b00100110000100001001111000011000;
		kmersSeqOne[14]= 32'b10011000010000100111100001100000;
		kmersSeqOne[15]= 32'b01100001000010011110000110000001;
		kmersSeqOne[16]= 32'b10000100001001111000011000000110;
		kmersSeqOne[17]= 32'b00010000100111100001100000011011;
		kmersSeqOne[18]= 32'b01000010011110000110000001101111;
		kmersSeqOne[19]= 32'b00001001111000011000000110111110;
		kmersSeqOne[20]= 32'b00100111100001100000011011111000;
		kmersSeqOne[21]= 32'b10011110000110000001101111100001;
		kmersSeqOne[22]= 32'b01111000011000000110111110000100;
		kmersSeqOne[23]= 32'b11100001100000011011111000010010;
		kmersSeqOne[24]= 32'b10000110000001101111100001001000;
		kmersSeqOne[25]= 32'b00011000000110111110000100100001;
		kmersSeqOne[26]= 32'b01100000011011111000010010000101;
		kmersSeqOne[27]= 32'b10000001101111100001001000010101;
		kmersSeqOne[28]= 32'b00000110111110000100100001010110;
		kmersSeqOne[29]= 32'b00011011111000010010000101011000;
		kmersSeqOne[30]= 32'b01101111100001001000010101100010;
		kmersSeqOne[31]= 32'b10111110000100100001010110001011;
		kmersSeqOne[32]= 32'b11111000010010000101011000101110;
		kmersSeqOne[33]= 32'b11100001001000010101100010111010;
		kmersSeqOne[34]= 32'b10000100100001010110001011101011;
		kmersSeqOne[35]= 32'b00010010000101011000101110101100;
		kmersSeqOne[36]= 32'b01001000010101100010111010110000;
		kmersSeqOne[37]= 32'b00100001010110001011101011000010;
		kmersSeqOne[38]= 32'b10000101011000101110101100001001;
		kmersSeqOne[39]= 32'b00010101100010111010110000100101;
		kmersSeqOne[40]= 32'b01010110001011101011000010010110;
		kmersSeqOne[41]= 32'b01011000101110101100001001011011;
		kmersSeqOne[42]= 32'b01100010111010110000100101101110;
		kmersSeqOne[43]= 32'b10001011101011000010010110111001;
		kmersSeqOne[44]= 32'b00101110101100001001011011100100;
		kmersSeqOne[45]= 32'b10111010110000100101101110010010;
		kmersSeqOne[46]= 32'b11101011000010010110111001001001;
		kmersSeqOne[47]= 32'b10101100001001011011100100100111;
		kmersSeqOne[48]= 32'b10110000100101101110010010011110;
		kmersSeqTwo[0]= 32'b10000111100001100111100010011111;
		kmersSeqTwo[1]= 32'b00011110000110011110001001111100;
		kmersSeqTwo[2]= 32'b01111000011001111000100111110010;
		kmersSeqTwo[3]= 32'b11100001100111100010011111001001;
		kmersSeqTwo[4]= 32'b10000110011110001001111100100111;
		kmersSeqTwo[5]= 32'b00011001111000100111110010011111;
		kmersSeqTwo[6]= 32'b01100111100010011111001001111111;
		kmersSeqTwo[7]= 32'b10011110001001111100100111111111;
		kmersSeqTwo[8]= 32'b01111000100111110010011111111111;
		kmersSeqTwo[9]= 32'b11100010011111001001111111111111;
		kmersSeqTwo[10]= 32'b10001001111100100111111111111111;
		kmersSeqTwo[11]= 32'b00100111110010011111111111111111;
		kmersSeqTwo[12]= 32'b10011111001001111111111111111111;
		kmersSeqTwo[13]= 32'b01111100100111111111111111111111;
		kmersSeqTwo[14]= 32'b11110010011111111111111111111111;
		kmersSeqTwo[15]= 32'b11001001111111111111111111111110;
		kmersSeqTwo[16]= 32'b00100111111111111111111111111000;
		kmersSeqTwo[17]= 32'b10011111111111111111111111100001;
		kmersSeqTwo[18]= 32'b01111111111111111111111110000110;
		kmersSeqTwo[19]= 32'b11111111111111111111111000011000;
		kmersSeqTwo[20]= 32'b11111111111111111111100001100001;
		kmersSeqTwo[21]= 32'b11111111111111111110000110000110;
		kmersSeqTwo[22]= 32'b11111111111111111000011000011000;
		kmersSeqTwo[23]= 32'b11111111111111100001100001100011;
		kmersSeqTwo[24]= 32'b11111111111110000110000110001110;
		kmersSeqTwo[25]= 32'b11111111111000011000011000111010;
		kmersSeqTwo[26]= 32'b11111111100001100001100011101001;
		kmersSeqTwo[27]= 32'b11111110000110000110001110100101;
		kmersSeqTwo[28]= 32'b11111000011000011000111010010110;
		kmersSeqTwo[29]= 32'b11100001100001100011101001011010;
		kmersSeqTwo[30]= 32'b10000110000110001110100101101000;
		kmersSeqTwo[31]= 32'b00011000011000111010010110100011;
		kmersSeqTwo[32]= 32'b01100001100011101001011010001111;
		kmersSeqTwo[33]= 32'b10000110001110100101101000111110;
		kmersSeqTwo[34]= 32'b00011000111010010110100011111011;
		kmersSeqTwo[35]= 32'b01100011101001011010001111101111;
		kmersSeqTwo[36]= 32'b10001110100101101000111110111111;
		kmersSeqTwo[37]= 32'b00111010010110100011111011111111;
		kmersSeqTwo[38]= 32'b11101001011010001111101111111111;
		kmersSeqTwo[39]= 32'b10100101101000111110111111111111;
		kmersSeqTwo[40]= 32'b10010110100011111011111111111111;
		kmersSeqTwo[41]= 32'b01011010001111101111111111111111;
		kmersSeqTwo[42]= 32'b01101000111110111111111111111111;
		kmersSeqTwo[43]= 32'b10100011111011111111111111111111;
		kmersSeqTwo[44]= 32'b10001111101111111111111111111100;
		kmersSeqTwo[45]= 32'b00111110111111111111111111110010;
		kmersSeqTwo[46]= 32'b11111011111111111111111111001001;
		kmersSeqTwo[47]= 32'b11101111111111111111111100100101;
		kmersSeqTwo[48]= 32'b10111111111111111111110010010110;
		#20 rstN = 0;
		randA =  10323 ;
		randB =  10091 ;
		#80
		randA =  2324 ;
		randB =  1 ;
		#80
		randA =  358771 ;
		randB =  233 ;
		#80
		randA =  409712 ;
		randB =  76423 ;
		#80
		randA =  94390 ;
		randB =  4232409 ;
		#80
		randA =  2229481 ;
		randB =  57554 ;
		#80
		randA =  123 ;
		randB =  2231130 ;
		#80
		randA =  1441 ;
		randB =  1091 ;
		#260
		rstN = 1;
		$stop;
		$finish;
	end
	
	
	
	endmodule
	