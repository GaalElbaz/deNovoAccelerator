module topDesgin_tbTwo();

	logic clk, rstN;
	logic [31:0] randA;
	logic [31:0] randB;
	logic unsigned [48:0][31:0] kmersSeqOne;
	logic unsigned [48:0][31:0] kmersSeqTwo;
	logic unsigned [4:0] jaccardSimilarity;
	
	topDesginModule myTopDesginTB(.clk(clk), .rstN(rstN), .randA(randA), .randB(randB), .kmersSeqOne(kmersSeqOne), .kmersSeqTwo(kmersSeqTwo), .jaccardSimilarity(jaccardSimilarity));
	
	always begin
		#40 clk = ~clk;
	end
	
	initial begin
		clk = 0;
		rstN = 1;
			kmersSeqOne[0]= 32'b11111111111111111111111111111111;
		kmersSeqOne[1]= 32'b11111111111111111111111111111111;
		kmersSeqOne[2]= 32'b11111111111111111111111111111111;
		kmersSeqOne[3]= 32'b11111111111111111111111111111111;
		kmersSeqOne[4]= 32'b11111111111111111111111111111111;
		kmersSeqOne[5]= 32'b11111111111111111111111111111111;
		kmersSeqOne[6]= 32'b11111111111111111111111111111111;
		kmersSeqOne[7]= 32'b11111111111111111111111111111111;
		kmersSeqOne[8]= 32'b11111111111111111111111111111111;
		kmersSeqOne[9]= 32'b11111111111111111111111111111111;
		kmersSeqOne[10]= 32'b11111111111111111111111111111111;
		kmersSeqOne[11]= 32'b11111111111111111111111111111111;
		kmersSeqOne[12]= 32'b11111111111111111111111111111111;
		kmersSeqOne[13]= 32'b11111111111111111111111111111111;
		kmersSeqOne[14]= 32'b11111111111111111111111111111111;
		kmersSeqOne[15]= 32'b11111111111111111111111111111111;
		kmersSeqOne[16]= 32'b11111111111111111111111111111111;
		kmersSeqOne[17]= 32'b11111111111111111111111111111111;
		kmersSeqOne[18]= 32'b11111111111111111111111111111111;
		kmersSeqOne[19]= 32'b11111111111111111111111111111111;
		kmersSeqOne[20]= 32'b11111111111111111111111111111111;
		kmersSeqOne[21]= 32'b11111111111111111111111111111111;
		kmersSeqOne[22]= 32'b11111111111111111111111111111111;
		kmersSeqOne[23]= 32'b11111111111111111111111111111111;
		kmersSeqOne[24]= 32'b11111111111111111111111111111111;
		kmersSeqOne[25]= 32'b11111111111111111111111111111111;
		kmersSeqOne[26]= 32'b11111111111111111111111111111111;
		kmersSeqOne[27]= 32'b11111111111111111111111111111111;
		kmersSeqOne[28]= 32'b11111111111111111111111111111111;
		kmersSeqOne[29]= 32'b11111111111111111111111111111111;
		kmersSeqOne[30]= 32'b11111111111111111111111111111111;
		kmersSeqOne[31]= 32'b11111111111111111111111111111111;
		kmersSeqOne[32]= 32'b11111111111111111111111111111111;
		kmersSeqOne[33]= 32'b11111111111111111111111111111111;
		kmersSeqOne[34]= 32'b11111111111111111111111111111111;
		kmersSeqOne[35]= 32'b11111111111111111111111111111111;
		kmersSeqOne[36]= 32'b11111111111111111111111111111111;
		kmersSeqOne[37]= 32'b11111111111111111111111111111111;
		kmersSeqOne[38]= 32'b11111111111111111111111111111111;
		kmersSeqOne[39]= 32'b11111111111111111111111111111111;
		kmersSeqOne[40]= 32'b11111111111111111111111111111111;
		kmersSeqOne[41]= 32'b11111111111111111111111111111111;
		kmersSeqOne[42]= 32'b11111111111111111111111111111111;
		kmersSeqOne[43]= 32'b11111111111111111111111111111111;
		kmersSeqOne[44]= 32'b11111111111111111111111111111111;
		kmersSeqOne[45]= 32'b11111111111111111111111111111111;
		kmersSeqOne[46]= 32'b11111111111111111111111111111111;
		kmersSeqOne[47]= 32'b11111111111111111111111111111111;
		kmersSeqOne[48]= 32'b11111111111111111111111111111111;
		kmersSeqTwo[0]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[1]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[2]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[3]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[4]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[5]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[6]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[7]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[8]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[9]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[10]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[11]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[12]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[13]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[14]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[15]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[16]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[17]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[18]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[19]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[20]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[21]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[22]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[23]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[24]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[25]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[26]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[27]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[28]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[29]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[30]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[31]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[32]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[33]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[34]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[35]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[36]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[37]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[38]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[39]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[40]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[41]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[42]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[43]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[44]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[45]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[46]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[47]= 32'b00000000000000000000000000000000;
		kmersSeqTwo[48]= 32'b00000000000000000000000000000000;
		#20 rstN = 0;
		randA =  10323 ;
		randB =  10091 ;
		#80
		randA =  2324 ;
		randB =  1 ;
		#80
		randA =  358771 ;
		randB =  233 ;
		#80
		randA =  409712 ;
		randB =  76423 ;
		#80
		randA =  94390 ;
		randB =  4232409 ;
		#80
		randA =  2229481 ;
		randB =  57554 ;
		#80
		randA =  123 ;
		randB =  2231130 ;
		#80
		randA =  1441 ;
		randB =  1091 ;
		#260
		rstN = 1;
		$stop;
		$finish;
	end
	
	
	
	endmodule
	
